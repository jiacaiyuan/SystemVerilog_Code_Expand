`define RID_WIDTH_NEST   100